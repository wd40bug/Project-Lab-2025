`timescale 1ns/1ps
module ClawServo_tb();
endmodule
